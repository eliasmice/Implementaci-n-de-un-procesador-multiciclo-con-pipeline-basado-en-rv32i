
// ALU

module alu(
input logic   [31:0] SrcA, 
input logic   [31:0] SrcB, 
input logic   [3:0]  ALUControl , 
output logic  [31:0] ALUResult, 
output logic         Zero, Sign);

logic [31:0] Sum;
logic Overflow;

assign Sum = SrcA + (ALUControl[0] ? ~SrcB : SrcB) + ALUControl[0];  // sub using 1's complement
assign Overflow = ~(ALUControl[0] ^ SrcB[31] ^ SrcA[31]) & (SrcA[31] ^ Sum[31]) & (~ALUControl[1]);

assign Zero = ~(|ALUResult);
assign Sign = ALUResult[31];

always_comb
		casex (ALUControl)
				4'b000x: ALUResult = Sum;				                  // sum or diff
				4'b0010: ALUResult = SrcA & SrcB;	                      // and
				4'b0011: ALUResult = SrcA | SrcB;	                      // or
				4'b0100: ALUResult = SrcA << SrcB;	                      // sll, slli
				4'b0101: ALUResult = {{30{1'b0}}, Overflow ^ Sum[31]};    //slt, slti
				4'b0110: ALUResult = SrcA ^ SrcB;                         // Xor
				4'b0111: ALUResult = SrcA >> SrcB;                        // shift logic
				4'b1000: ALUResult = ($unsigned(SrcA) < $unsigned(SrcB)); //sltu, stlui
				4'b1111: ALUResult = SrcA >>> SrcB;                       //shift arithmetic
				default: ALUResult = 32'bx;
		endcase
endmodule